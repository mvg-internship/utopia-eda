module NAND(A, B, Y);
input A, B;
output Y = ~(A & B);
endmodule




