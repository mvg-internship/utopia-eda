module A(a,c);
input a;
output c;
not n1(c,b);
endmodule

