/*Incorrect order of signals in not gates*/

module s344(GND,VDD,CK,A0,A1,A2,A3,B0,B1,B2,B3,CNTVCO2,CNTVCON2,P0,P1,P2,P3,P4,
  P5,P6,P7,READY,START);
input GND,VDD,CK,START,B0,B1,B2,B3,A0,A1,A2,A3;
output P4,P5,P6,P7,P0,P1,P2,P3,CNTVCON2,CNTVCO2,READY;

  wire CT2,CNTVG3VD,CT1,CNTVG2VD,CT0,CNTVG1VD,ACVQN3,ACVG4VD1,ACVQN2,ACVG3VD1,
    ACVQN1,ACVG2VD1,ACVQN0,ACVG1VD1,MRVQN3,MRVG4VD,MRVQN2,MRVG3VD,MRVQN1,
    MRVG2VD,MRVQN0,MRVG1VD,AX3,AM3,AX2,AM2,AX1,AM1,AX0,AM0,CNTVG3VQN,CNTVG2VQN,
    CNTVG1VQN,CNTVCON0,CT1N,ACVPCN,CNTVCO0,AMVS0N,IINIIT,READYN,BMVS0N,
    AMVG5VS0P,AMVG4VS0P,AMVG3VS0P,AMVG2VS0P,AD0,AD0N,AD1,AD1N,AD2,AD2N,AD3,
    AD3N,CNTVG3VD1,CNTVCON1,CNTVG1VD1,BMVG5VS0P,BMVG4VS0P,BMVG3VS0P,BMVG2VS0P,
    SMVS0N,ADSH,MRVSHLDN,ADDVC1,ADDVG1VCN,SMVG5VS0P,SMVG4VS0P,SMVG3VS0P,
    SMVG2VS0P,CNTVG1VZ,CNTVG1VZ1,AMVG5VX,AMVG4VX,AMVG3VX,AMVG2VX,S0,ADDVG1VP,
    BM3,BMVG5VX,BM2,BMVG4VX,BM1,BMVG3VX,BM0,BMVG2VX,ADDVC2,ADDVG2VCN,S1,
    ADDVG2VSN,ADDVC3,ADDVG3VCN,S2,ADDVG3VSN,SM0,SMVG2VX,CO,ADDVG4VCN,S3,
    ADDVG4VSN,SM1,SMVG3VX,SM3,SMVG5VX,SM2,SMVG4VX,AMVG5VG1VAD1NF,
    AMVG4VG1VAD1NF,AMVG3VG1VAD1NF,AMVG2VG1VAD1NF,BMVG5VG1VAD1NF,BMVG4VG1VAD1NF,
    BMVG3VG1VAD1NF,BMVG2VG1VAD1NF,AMVG5VG1VAD2NF,AMVG4VG1VAD2NF,AMVG3VG1VAD2NF,
    AMVG2VG1VAD2NF,ADDVG2VCNVAD1NF,ADDVG3VCNVAD1NF,ADDVG4VCNVAD1NF,
    MRVG3VDVAD1NF,MRVG2VDVAD1NF,MRVG1VDVAD1NF,BMVG5VG1VAD2NF,BMVG4VG1VAD2NF,
    BMVG3VG1VAD2NF,BMVG2VG1VAD2NF,SMVG5VG1VAD1NF,SMVG4VG1VAD1NF,SMVG3VG1VAD1NF,
    SMVG2VG1VAD1NF,ADDVG2VCNVAD4NF,ADDVG2VCNVAD2NF,ADDVG2VCNVOR1NF,
    MRVG4VDVAD1NF,MRVG4VDVAD2NF,MRVG3VDVAD2NF,MRVG2VDVAD2NF,MRVG1VDVAD2NF,
    ADDVG2VCNVAD3NF,ADDVG2VCNVOR2NF,ADDVG3VCNVAD4NF,ADDVG3VCNVAD2NF,
    ADDVG3VCNVOR1NF,ADDVG3VCNVAD3NF,ADDVG3VCNVOR2NF,SMVG2VG1VAD2NF,
    ADDVG4VCNVAD4NF,ADDVG4VCNVAD2NF,ADDVG4VCNVOR1NF,ADDVG4VCNVAD3NF,
    ADDVG4VCNVOR2NF,SMVG3VG1VAD2NF,SMVG5VG1VAD2NF,SMVG4VG1VAD2NF,
    ADDVG1VPVOR1NF,CNTVG3VG2VOR1NF,CNTVG2VG2VOR1NF,CNTVG2VD1,CNTVCO1,CNTVG3VZ1,
    CNTVG2VZ1,CNTVG3VZ,CNTVG2VZ;

  dff DFF_0(CK,CT2,CNTVG3VD);
  dff DFF_1(CK,CT1,CNTVG2VD);
  dff DFF_2(CK,CT0,CNTVG1VD);
  dff DFF_3(CK,ACVQN3,ACVG4VD1);
  dff DFF_4(CK,ACVQN2,ACVG3VD1);
  dff DFF_5(CK,ACVQN1,ACVG2VD1);
  dff DFF_6(CK,ACVQN0,ACVG1VD1);
  dff DFF_7(CK,MRVQN3,MRVG4VD);
  dff DFF_8(CK,MRVQN2,MRVG3VD);
  dff DFF_9(CK,MRVQN1,MRVG2VD);
  dff DFF_10(CK,MRVQN0,MRVG1VD);
  dff DFF_11(CK,AX3,AM3);
  dff DFF_12(CK,AX2,AM2);
  dff DFF_13(CK,AX1,AM1);
  dff DFF_14(CK,AX0,AM0);
  not NOT_0(CNTVG3VQN,CT2);
  not NOT_1(CNTVG2VQN,CT1);
  not NOT_2(CNTVG1VQN,CT0);
  not NOT_3(P7,ACVQN3);
  not NOT_4(P6,ACVQN2);
  not NOT_5(P5,ACVQN1);
  not NOT_6(P4,ACVQN0);
  not NOT_7(P3,MRVQN3);
  not NOT_8(P2,MRVQN2);
  not NOT_9(P1,MRVQN1);
  not NOT_10(P0,MRVQN0);
  not NOT_11(CNTVCON0,CT0);
  not NOT_12(CT1N,CT1);
  not NOT_13(ACVPCN,START);
  not NOT_14(CNTVCO0,CNTVG1VQN);
  not NOT_15(AMVS0N,IINIIT);
  not NOT_16(READY,READYN);
  not NOT_17(BMVS0N,READYN);
  not NOT_18(AMVG5VS0P,AMVS0N);
  not NOT_19(AMVG4VS0P,AMVS0N);
  not NOT_20(AMVG3VS0P,AMVS0N);
  not NOT_21(AMVG2VS0P,AMVS0N);
  not NOT_22(AD0,AD0N);
  not NOT_23(AD1,AD1N);
  not NOT_24(AD2,AD2N);
  not NOT_25(AD3,AD3N);
  not NOT_26(CNTVG3VD1,CNTVCON1);
  not NOT_27(CNTVG1VD1,READY);
  not NOT_28(BMVG5VS0P,BMVS0N);
  not NOT_29(BMVG4VS0P,BMVS0N);
  not NOT_30(BMVG3VS0P,BMVS0N);
  not NOT_31(BMVG2VS0P,BMVS0N);
  not NOT_32(SMVS0N,ADSH);
  not NOT_33(MRVSHLDN,ADSH);
  not NOT_34(ADDVC1,ADDVG1VCN);
  not NOT_35(SMVG5VS0P,SMVS0N);
  not NOT_36(SMVG4VS0P,SMVS0N);
  not NOT_37(SMVG3VS0P,SMVS0N);
  not NOT_38(SMVG2VS0P,SMVS0N);
  not NOT_39(CNTVG1VZ,CNTVG1VZ1);
  not NOT_40(AM3,AMVG5VX);
  not NOT_41(AM2,AMVG4VX);
  not NOT_42(AM1,AMVG3VX);
  not NOT_43(AM0,AMVG2VX);
  not NOT_44(S0,ADDVG1VP);
  not NOT_45(BM3,BMVG5VX);
  not NOT_46(BM2,BMVG4VX);
  not NOT_47(BM1,BMVG3VX);
  not NOT_48(BM0,BMVG2VX);
  not NOT_49(ADDVC2,ADDVG2VCN);
  not NOT_50(S1,ADDVG2VSN);
  not NOT_51(ADDVC3,ADDVG3VCN);
  not NOT_52(S2,ADDVG3VSN);
  not NOT_53(SM0,SMVG2VX);
  not NOT_54(CO,ADDVG4VCN);
  not NOT_55(S3,ADDVG4VSN);
  not NOT_56(SM1,SMVG3VX);
  not NOT_57(SM3,SMVG5VX);
  not NOT_58(SM2,SMVG4VX);
  and AND2_0(AMVG5VG1VAD1NF,AMVS0N,AX3);
  and AND2_1(AMVG4VG1VAD1NF,AMVS0N,AX2);
  and AND2_2(AMVG3VG1VAD1NF,AMVS0N,AX1);
  and AND2_3(AMVG2VG1VAD1NF,AMVS0N,AX0);
  and AND2_4(BMVG5VG1VAD1NF,BMVS0N,P3);
  and AND2_5(BMVG4VG1VAD1NF,BMVS0N,P2);
  and AND2_6(BMVG3VG1VAD1NF,BMVS0N,P1);
  and AND2_7(BMVG2VG1VAD1NF,BMVS0N,P0);
  and AND2_8(AMVG5VG1VAD2NF,AMVG5VS0P,A3);
  and AND2_9(AMVG4VG1VAD2NF,AMVG4VS0P,A2);
  and AND2_10(AMVG3VG1VAD2NF,AMVG3VS0P,A1);
  and AND2_11(AMVG2VG1VAD2NF,AMVG2VS0P,A0);
  and AND2_12(ADDVG2VCNVAD1NF,AD1,P5);
  and AND2_13(ADDVG3VCNVAD1NF,AD2,P6);
  and AND2_14(ADDVG4VCNVAD1NF,AD3,P7);
  and AND2_15(MRVG3VDVAD1NF,ADSH,P3);
  and AND2_16(MRVG2VDVAD1NF,ADSH,P2);
  and AND2_17(MRVG1VDVAD1NF,ADSH,P1);
  and AND2_18(BMVG5VG1VAD2NF,BMVG5VS0P,B3);
  and AND2_19(BMVG4VG1VAD2NF,BMVG4VS0P,B2);
  and AND2_20(BMVG3VG1VAD2NF,BMVG3VS0P,B1);
  and AND2_21(BMVG2VG1VAD2NF,BMVG2VS0P,B0);
  and AND2_22(SMVG5VG1VAD1NF,SMVS0N,P7);
  and AND2_23(SMVG4VG1VAD1NF,SMVS0N,P6);
  and AND2_24(SMVG3VG1VAD1NF,SMVS0N,P5);
  and AND2_25(SMVG2VG1VAD1NF,SMVS0N,P4);
  and AND3_0(ADDVG2VCNVAD4NF,ADDVC1,AD1,P5);
  and AND2_26(ADDVG2VCNVAD2NF,ADDVC1,ADDVG2VCNVOR1NF);
  and AND2_27(MRVG4VDVAD1NF,ADSH,S0);
  and AND2_28(MRVG4VDVAD2NF,MRVSHLDN,BM3);
  and AND2_29(MRVG3VDVAD2NF,MRVSHLDN,BM2);
  and AND2_30(MRVG2VDVAD2NF,MRVSHLDN,BM1);
  and AND2_31(MRVG1VDVAD2NF,MRVSHLDN,BM0);
  and AND2_32(ADDVG2VCNVAD3NF,ADDVG2VCNVOR2NF,ADDVG2VCN);
  and AND3_1(ADDVG3VCNVAD4NF,ADDVC2,AD2,P6);
  and AND2_33(ADDVG3VCNVAD2NF,ADDVC2,ADDVG3VCNVOR1NF);
  and AND2_34(ADDVG3VCNVAD3NF,ADDVG3VCNVOR2NF,ADDVG3VCN);
  and AND2_35(SMVG2VG1VAD2NF,SMVG2VS0P,S1);
  and AND3_2(ADDVG4VCNVAD4NF,ADDVC3,AD3,P7);
  and AND2_36(ADDVG4VCNVAD2NF,ADDVC3,ADDVG4VCNVOR1NF);
  and AND2_37(ADDVG4VCNVAD3NF,ADDVG4VCNVOR2NF,ADDVG4VCN);
  and AND2_38(SMVG3VG1VAD2NF,SMVG3VS0P,S2);
  and AND2_39(SMVG5VG1VAD2NF,SMVG5VS0P,CO);
  and AND2_40(SMVG4VG1VAD2NF,SMVG4VS0P,S3);
  or OR2_0(ADDVG1VPVOR1NF,AD0,P4);
  or OR2_1(ADDVG2VCNVOR1NF,AD1,P5);
  or OR2_2(ADDVG3VCNVOR1NF,AD2,P6);
  or OR2_3(ADDVG4VCNVOR1NF,AD3,P7);
  or OR2_4(CNTVG3VG2VOR1NF,CT2,CNTVG3VD1);
  or OR2_5(CNTVG2VG2VOR1NF,CT1,CNTVG2VD1);
  or OR3_0(ADDVG2VCNVOR2NF,ADDVC1,AD1,P5);
  or OR3_1(ADDVG3VCNVOR2NF,ADDVC2,AD2,P6);
  or OR3_2(ADDVG4VCNVOR2NF,ADDVC3,AD3,P7);
  nand NAND3_0(READYN,CT0,CT1N,CT2);
  nand NAND2_0(AD0N,P0,AX0);
  nand NAND2_1(AD1N,P0,AX1);
  nand NAND2_2(AD2N,P0,AX2);
  nand NAND2_3(AD3N,P0,AX3);
  nand NAND2_4(CNTVCON1,CT1,CNTVCO0);
  nand NAND2_5(CNTVCON2,CT2,CNTVCO1);
  nand NAND2_6(ADDVG1VCN,AD0,P4);
  nand NAND2_7(CNTVG3VZ1,CT2,CNTVG3VD1);
  nand NAND2_8(CNTVG2VZ1,CT1,CNTVG2VD1);
  nand NAND2_9(CNTVG1VZ1,CT0,CNTVG1VD1);
  nand NAND2_10(ADDVG1VP,ADDVG1VPVOR1NF,ADDVG1VCN);
  nand NAND2_11(CNTVG3VZ,CNTVG3VG2VOR1NF,CNTVG3VZ1);
  nand NAND2_12(CNTVG2VZ,CNTVG2VG2VOR1NF,CNTVG2VZ1);
  nand NAND2_13(ACVG1VD1,ACVPCN,SM0);
  nand NAND2_14(ACVG2VD1,ACVPCN,SM1);
  nand NAND2_15(ACVG4VD1,ACVPCN,SM3);
  nand NAND2_16(ACVG3VD1,ACVPCN,SM2);
  nor NOR3_0(IINIIT,CT0,CT1,CT2);
  nor NOR2_0(CNTVCO1,CNTVG2VQN,CNTVCON0);
  nor NOR2_1(CNTVCO2,CNTVG3VQN,CNTVCON1);
  nor NOR2_2(ADSH,READY,IINIIT);
  nor NOR2_3(CNTVG2VD1,READY,CNTVCON0);
  nor NOR2_4(AMVG5VX,AMVG5VG1VAD2NF,AMVG5VG1VAD1NF);
  nor NOR2_5(AMVG4VX,AMVG4VG1VAD2NF,AMVG4VG1VAD1NF);
  nor NOR2_6(AMVG3VX,AMVG3VG1VAD2NF,AMVG3VG1VAD1NF);
  nor NOR2_7(AMVG2VX,AMVG2VG1VAD2NF,AMVG2VG1VAD1NF);
  nor NOR2_8(BMVG5VX,BMVG5VG1VAD2NF,BMVG5VG1VAD1NF);
  nor NOR2_9(BMVG4VX,BMVG4VG1VAD2NF,BMVG4VG1VAD1NF);
  nor NOR2_10(BMVG3VX,BMVG3VG1VAD2NF,BMVG3VG1VAD1NF);
  nor NOR2_11(BMVG2VX,BMVG2VG1VAD2NF,BMVG2VG1VAD1NF);
  nor NOR2_12(CNTVG3VD,CNTVG3VZ,START);
  nor NOR2_13(CNTVG2VD,CNTVG2VZ,START);
  nor NOR2_14(CNTVG1VD,CNTVG1VZ,START);
  nor NOR2_15(ADDVG2VCN,ADDVG2VCNVAD2NF,ADDVG2VCNVAD1NF);
  nor NOR2_16(MRVG4VD,MRVG4VDVAD2NF,MRVG4VDVAD1NF);
  nor NOR2_17(MRVG3VD,MRVG3VDVAD2NF,MRVG3VDVAD1NF);
  nor NOR2_18(MRVG2VD,MRVG2VDVAD2NF,MRVG2VDVAD1NF);
  nor NOR2_19(MRVG1VD,MRVG1VDVAD2NF,MRVG1VDVAD1NF);
  nor NOR2_20(ADDVG2VSN,ADDVG2VCNVAD4NF,ADDVG2VCNVAD3NF);
  nor NOR2_21(ADDVG3VCN,ADDVG3VCNVAD2NF,ADDVG3VCNVAD1NF);
  nor NOR2_22(ADDVG3VSN,ADDVG3VCNVAD4NF,ADDVG3VCNVAD3NF);
  nor NOR2_23(SMVG2VX,SMVG2VG1VAD2NF,SMVG2VG1VAD1NF);
  nor NOR2_24(ADDVG4VCN,ADDVG4VCNVAD2NF,ADDVG4VCNVAD1NF);
  nor NOR2_25(ADDVG4VSN,ADDVG4VCNVAD4NF,ADDVG4VCNVAD3NF);
  nor NOR2_26(SMVG3VX,SMVG3VG1VAD2NF,SMVG3VG1VAD1NF);
  nor NOR2_27(SMVG5VX,SMVG5VG1VAD2NF,SMVG5VG1VAD1NF);
  nor NOR2_28(SMVG4VX,SMVG4VG1VAD2NF,SMVG4VG1VAD1NF);

endmodule