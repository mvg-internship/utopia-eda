module A(a,b);
input a;
output b;
not n1(b,a);
endmodule