module A(a,b,c);
input a,b;
output c;
xor x1(c,a,b);
endmodule