module A(a,b,c);
input a,b;
output c;
xnor xnr1(c,a,b);
endmodule