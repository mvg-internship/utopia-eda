module A(a,b,c);
input a,b;
output c;
nor nr1(c,a,b);
endmodule