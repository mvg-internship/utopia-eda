module orGate(cOut, x0, x1);
  input x0, x1, x2;
  output cOut;
  wire cOut;

  or g4 (cOut, x0, x1);
endmodule

