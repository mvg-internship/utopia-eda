module A(a,b,c);
input a,b;
output c;
or o1(c,a,b);
endmodule