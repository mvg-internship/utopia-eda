module SUM(A, C, Y);
input A,C;
output Y = A+C;
endmodule
