module SUM(A, C, Y);
input A,C;
output Y = A+C;
endmodule

module DEC(A,C,Y);
input A,C;
output Y = A-C;
endmodule
