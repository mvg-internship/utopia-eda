module A(a,a,b,c);
input a,b;
output c;
dff d1(a,c,b);
endmodule