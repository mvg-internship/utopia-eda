module A(a,b,c);
input a,b;
output c;
nand nd1(c,a,b);
endmodule